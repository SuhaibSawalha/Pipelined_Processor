module testbech ();
							
	
endmodule