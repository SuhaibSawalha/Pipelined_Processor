module add (
    input [15:0] a,
    output [15:0] sum
);

    assign sum = a + ;

endmodule
